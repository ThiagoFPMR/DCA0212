library verilog;
use verilog.vl_types.all;
entity FlipFlopD4BitRegister_vlg_vec_tst is
end FlipFlopD4BitRegister_vlg_vec_tst;
