library verilog;
use verilog.vl_types.all;
entity MagnitudeComparator4Bit_vlg_vec_tst is
end MagnitudeComparator4Bit_vlg_vec_tst;
