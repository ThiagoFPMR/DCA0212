library verilog;
use verilog.vl_types.all;
entity MagnitudeComparator1Bit_vlg_vec_tst is
end MagnitudeComparator1Bit_vlg_vec_tst;
