library verilog;
use verilog.vl_types.all;
entity LatchD4BitRegister_vlg_vec_tst is
end LatchD4BitRegister_vlg_vec_tst;
