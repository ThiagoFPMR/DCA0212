library verilog;
use verilog.vl_types.all;
entity MagnitudeComparator8Bit_vlg_vec_tst is
end MagnitudeComparator8Bit_vlg_vec_tst;
